module main;
   initial $s1Assembler("try.txt");
endmodule
