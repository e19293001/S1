module main;
   initial $s1Assembler("tst/test_parser_pattern0004.txt");
endmodule
